// hps.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module hps (
		output wire         capture_clk_clk,               //      capture_clk.clk
		output wire         capture_clk_div8_clk,          // capture_clk_div8.clk
		input  wire         clk_clk,                       //              clk.clk
		input  wire [26:0]  f2h_sdram0_data_address,       //  f2h_sdram0_data.address
		input  wire [7:0]   f2h_sdram0_data_burstcount,    //                 .burstcount
		output wire         f2h_sdram0_data_waitrequest,   //                 .waitrequest
		output wire [255:0] f2h_sdram0_data_readdata,      //                 .readdata
		output wire         f2h_sdram0_data_readdatavalid, //                 .readdatavalid
		input  wire         f2h_sdram0_data_read,          //                 .read
		input  wire [255:0] f2h_sdram0_data_writedata,     //                 .writedata
		input  wire [31:0]  f2h_sdram0_data_byteenable,    //                 .byteenable
		input  wire         f2h_sdram0_data_write,         //                 .write
		input  wire         h2f_lw_waitrequest,            //           h2f_lw.waitrequest
		input  wire [31:0]  h2f_lw_readdata,               //                 .readdata
		input  wire         h2f_lw_readdatavalid,          //                 .readdatavalid
		output wire [0:0]   h2f_lw_burstcount,             //                 .burstcount
		output wire [31:0]  h2f_lw_writedata,              //                 .writedata
		output wire [3:0]   h2f_lw_address,                //                 .address
		output wire         h2f_lw_write,                  //                 .write
		output wire         h2f_lw_read,                   //                 .read
		output wire [3:0]   h2f_lw_byteenable,             //                 .byteenable
		output wire         h2f_lw_debugaccess,            //                 .debugaccess
		output wire         mem_clk_clk,                   //          mem_clk.clk
		output wire [14:0]  memory_mem_a,                  //           memory.mem_a
		output wire [2:0]   memory_mem_ba,                 //                 .mem_ba
		output wire         memory_mem_ck,                 //                 .mem_ck
		output wire         memory_mem_ck_n,               //                 .mem_ck_n
		output wire         memory_mem_cke,                //                 .mem_cke
		output wire         memory_mem_cs_n,               //                 .mem_cs_n
		output wire         memory_mem_ras_n,              //                 .mem_ras_n
		output wire         memory_mem_cas_n,              //                 .mem_cas_n
		output wire         memory_mem_we_n,               //                 .mem_we_n
		output wire         memory_mem_reset_n,            //                 .mem_reset_n
		inout  wire [31:0]  memory_mem_dq,                 //                 .mem_dq
		inout  wire [3:0]   memory_mem_dqs,                //                 .mem_dqs
		inout  wire [3:0]   memory_mem_dqs_n,              //                 .mem_dqs_n
		output wire         memory_mem_odt,                //                 .mem_odt
		output wire [3:0]   memory_mem_dm,                 //                 .mem_dm
		input  wire         memory_oct_rzqin               //                 .oct_rzqin
	);

	wire  [63:0] pll_capture_reconfig_from_pll_reconfig_from_pll;                // pll_capture:reconfig_from_pll -> pll_reconfig_0:reconfig_from_pll
	wire  [63:0] pll_reconfig_0_reconfig_to_pll_reconfig_to_pll;                 // pll_reconfig_0:reconfig_to_pll -> pll_capture:reconfig_to_pll
	wire         hps_0_h2f_reset_reset;                                          // hps_0:h2f_rst_n -> [pll_capture:rst, pll_mem:rst, rst_controller:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                  // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                  // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                 // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                  // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                    // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                 // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                 // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                 // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                 // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                  // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                   // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                 // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                 // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                 // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                 // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                 // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                  // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                   // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                 // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata;    // pll_reconfig_0:mgmt_readdata -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest; // pll_reconfig_0:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_address -> pll_reconfig_0:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_read -> pll_reconfig_0:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_write -> pll_reconfig_0:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_writedata -> pll_reconfig_0:mgmt_writedata
	wire  [31:0] mm_interconnect_0_mm_bridge_h2f_lw_s0_readdata;                 // mm_bridge_h2f_lw:s0_readdata -> mm_interconnect_0:mm_bridge_h2f_lw_s0_readdata
	wire         mm_interconnect_0_mm_bridge_h2f_lw_s0_waitrequest;              // mm_bridge_h2f_lw:s0_waitrequest -> mm_interconnect_0:mm_bridge_h2f_lw_s0_waitrequest
	wire         mm_interconnect_0_mm_bridge_h2f_lw_s0_debugaccess;              // mm_interconnect_0:mm_bridge_h2f_lw_s0_debugaccess -> mm_bridge_h2f_lw:s0_debugaccess
	wire   [3:0] mm_interconnect_0_mm_bridge_h2f_lw_s0_address;                  // mm_interconnect_0:mm_bridge_h2f_lw_s0_address -> mm_bridge_h2f_lw:s0_address
	wire         mm_interconnect_0_mm_bridge_h2f_lw_s0_read;                     // mm_interconnect_0:mm_bridge_h2f_lw_s0_read -> mm_bridge_h2f_lw:s0_read
	wire   [3:0] mm_interconnect_0_mm_bridge_h2f_lw_s0_byteenable;               // mm_interconnect_0:mm_bridge_h2f_lw_s0_byteenable -> mm_bridge_h2f_lw:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_h2f_lw_s0_readdatavalid;            // mm_bridge_h2f_lw:s0_readdatavalid -> mm_interconnect_0:mm_bridge_h2f_lw_s0_readdatavalid
	wire         mm_interconnect_0_mm_bridge_h2f_lw_s0_write;                    // mm_interconnect_0:mm_bridge_h2f_lw_s0_write -> mm_bridge_h2f_lw:s0_write
	wire  [31:0] mm_interconnect_0_mm_bridge_h2f_lw_s0_writedata;                // mm_interconnect_0:mm_bridge_h2f_lw_s0_writedata -> mm_bridge_h2f_lw:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_bridge_h2f_lw_s0_burstcount;               // mm_interconnect_0:mm_bridge_h2f_lw_s0_burstcount -> mm_bridge_h2f_lw:s0_burstcount
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [mm_bridge_h2f_lw:reset, mm_interconnect_0:pll_reconfig_0_mgmt_reset_reset_bridge_in_reset_reset, pll_reconfig_0:mgmt_reset]

	hps_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.f2h_sdram0_clk           (mem_clk_clk),                     //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (f2h_sdram0_data_address),         //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (f2h_sdram0_data_burstcount),      //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (f2h_sdram0_data_waitrequest),     //                  .waitrequest
		.f2h_sdram0_READDATA      (f2h_sdram0_data_readdata),        //                  .readdata
		.f2h_sdram0_READDATAVALID (f2h_sdram0_data_readdatavalid),   //                  .readdatavalid
		.f2h_sdram0_READ          (f2h_sdram0_data_read),            //                  .read
		.f2h_sdram0_WRITEDATA     (f2h_sdram0_data_writedata),       //                  .writedata
		.f2h_sdram0_BYTEENABLE    (f2h_sdram0_data_byteenable),      //                  .byteenable
		.f2h_sdram0_WRITE         (f2h_sdram0_data_write),           //                  .write
		.h2f_axi_clk              (mem_clk_clk),                     //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                //                  .awaddr
		.h2f_AWLEN                (),                                //                  .awlen
		.h2f_AWSIZE               (),                                //                  .awsize
		.h2f_AWBURST              (),                                //                  .awburst
		.h2f_AWLOCK               (),                                //                  .awlock
		.h2f_AWCACHE              (),                                //                  .awcache
		.h2f_AWPROT               (),                                //                  .awprot
		.h2f_AWVALID              (),                                //                  .awvalid
		.h2f_AWREADY              (),                                //                  .awready
		.h2f_WID                  (),                                //                  .wid
		.h2f_WDATA                (),                                //                  .wdata
		.h2f_WSTRB                (),                                //                  .wstrb
		.h2f_WLAST                (),                                //                  .wlast
		.h2f_WVALID               (),                                //                  .wvalid
		.h2f_WREADY               (),                                //                  .wready
		.h2f_BID                  (),                                //                  .bid
		.h2f_BRESP                (),                                //                  .bresp
		.h2f_BVALID               (),                                //                  .bvalid
		.h2f_BREADY               (),                                //                  .bready
		.h2f_ARID                 (),                                //                  .arid
		.h2f_ARADDR               (),                                //                  .araddr
		.h2f_ARLEN                (),                                //                  .arlen
		.h2f_ARSIZE               (),                                //                  .arsize
		.h2f_ARBURST              (),                                //                  .arburst
		.h2f_ARLOCK               (),                                //                  .arlock
		.h2f_ARCACHE              (),                                //                  .arcache
		.h2f_ARPROT               (),                                //                  .arprot
		.h2f_ARVALID              (),                                //                  .arvalid
		.h2f_ARREADY              (),                                //                  .arready
		.h2f_RID                  (),                                //                  .rid
		.h2f_RDATA                (),                                //                  .rdata
		.h2f_RRESP                (),                                //                  .rresp
		.h2f_RLAST                (),                                //                  .rlast
		.h2f_RVALID               (),                                //                  .rvalid
		.h2f_RREADY               (),                                //                  .rready
		.h2f_lw_axi_clk           (mem_clk_clk),                     //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (4),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_h2f_lw (
		.clk              (mem_clk_clk),                                         //   clk.clk
		.reset            (rst_controller_reset_out_reset),                      // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_h2f_lw_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_h2f_lw_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_h2f_lw_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_h2f_lw_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_h2f_lw_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_h2f_lw_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_h2f_lw_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_h2f_lw_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_h2f_lw_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_h2f_lw_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (h2f_lw_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (h2f_lw_readdata),                                     //      .readdata
		.m0_readdatavalid (h2f_lw_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (h2f_lw_burstcount),                                   //      .burstcount
		.m0_writedata     (h2f_lw_writedata),                                    //      .writedata
		.m0_address       (h2f_lw_address),                                      //      .address
		.m0_write         (h2f_lw_write),                                        //      .write
		.m0_read          (h2f_lw_read),                                         //      .read
		.m0_byteenable    (h2f_lw_byteenable),                                   //      .byteenable
		.m0_debugaccess   (h2f_lw_debugaccess),                                  //      .debugaccess
		.s0_response      (),                                                    // (terminated)
		.m0_response      (2'b00)                                                // (terminated)
	);

	hps_pll_capture pll_capture (
		.refclk            (clk_clk),                                         //            refclk.clk
		.rst               (~hps_0_h2f_reset_reset),                          //             reset.reset
		.outclk_0          (capture_clk_clk),                                 //           outclk0.clk
		.outclk_1          (capture_clk_div8_clk),                            //           outclk1.clk
		.locked            (),                                                //            locked.export
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll),  //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_capture_reconfig_from_pll_reconfig_from_pll)  // reconfig_from_pll.reconfig_from_pll
	);

	hps_pll_mem pll_mem (
		.refclk   (clk_clk),                //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset), //   reset.reset
		.outclk_0 (mem_clk_clk),            // outclk0.clk
		.locked   ()                        //  locked.export
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_0 (
		.mgmt_clk          (mem_clk_clk),                                                    //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_reset_out_reset),                                 //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_capture_reconfig_from_pll_reconfig_from_pll),                // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	hps_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                          (hps_0_h2f_lw_axi_master_awid),                                   //                         hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                        (hps_0_h2f_lw_axi_master_awaddr),                                 //                                                .awaddr
		.hps_0_h2f_lw_axi_master_awlen                         (hps_0_h2f_lw_axi_master_awlen),                                  //                                                .awlen
		.hps_0_h2f_lw_axi_master_awsize                        (hps_0_h2f_lw_axi_master_awsize),                                 //                                                .awsize
		.hps_0_h2f_lw_axi_master_awburst                       (hps_0_h2f_lw_axi_master_awburst),                                //                                                .awburst
		.hps_0_h2f_lw_axi_master_awlock                        (hps_0_h2f_lw_axi_master_awlock),                                 //                                                .awlock
		.hps_0_h2f_lw_axi_master_awcache                       (hps_0_h2f_lw_axi_master_awcache),                                //                                                .awcache
		.hps_0_h2f_lw_axi_master_awprot                        (hps_0_h2f_lw_axi_master_awprot),                                 //                                                .awprot
		.hps_0_h2f_lw_axi_master_awvalid                       (hps_0_h2f_lw_axi_master_awvalid),                                //                                                .awvalid
		.hps_0_h2f_lw_axi_master_awready                       (hps_0_h2f_lw_axi_master_awready),                                //                                                .awready
		.hps_0_h2f_lw_axi_master_wid                           (hps_0_h2f_lw_axi_master_wid),                                    //                                                .wid
		.hps_0_h2f_lw_axi_master_wdata                         (hps_0_h2f_lw_axi_master_wdata),                                  //                                                .wdata
		.hps_0_h2f_lw_axi_master_wstrb                         (hps_0_h2f_lw_axi_master_wstrb),                                  //                                                .wstrb
		.hps_0_h2f_lw_axi_master_wlast                         (hps_0_h2f_lw_axi_master_wlast),                                  //                                                .wlast
		.hps_0_h2f_lw_axi_master_wvalid                        (hps_0_h2f_lw_axi_master_wvalid),                                 //                                                .wvalid
		.hps_0_h2f_lw_axi_master_wready                        (hps_0_h2f_lw_axi_master_wready),                                 //                                                .wready
		.hps_0_h2f_lw_axi_master_bid                           (hps_0_h2f_lw_axi_master_bid),                                    //                                                .bid
		.hps_0_h2f_lw_axi_master_bresp                         (hps_0_h2f_lw_axi_master_bresp),                                  //                                                .bresp
		.hps_0_h2f_lw_axi_master_bvalid                        (hps_0_h2f_lw_axi_master_bvalid),                                 //                                                .bvalid
		.hps_0_h2f_lw_axi_master_bready                        (hps_0_h2f_lw_axi_master_bready),                                 //                                                .bready
		.hps_0_h2f_lw_axi_master_arid                          (hps_0_h2f_lw_axi_master_arid),                                   //                                                .arid
		.hps_0_h2f_lw_axi_master_araddr                        (hps_0_h2f_lw_axi_master_araddr),                                 //                                                .araddr
		.hps_0_h2f_lw_axi_master_arlen                         (hps_0_h2f_lw_axi_master_arlen),                                  //                                                .arlen
		.hps_0_h2f_lw_axi_master_arsize                        (hps_0_h2f_lw_axi_master_arsize),                                 //                                                .arsize
		.hps_0_h2f_lw_axi_master_arburst                       (hps_0_h2f_lw_axi_master_arburst),                                //                                                .arburst
		.hps_0_h2f_lw_axi_master_arlock                        (hps_0_h2f_lw_axi_master_arlock),                                 //                                                .arlock
		.hps_0_h2f_lw_axi_master_arcache                       (hps_0_h2f_lw_axi_master_arcache),                                //                                                .arcache
		.hps_0_h2f_lw_axi_master_arprot                        (hps_0_h2f_lw_axi_master_arprot),                                 //                                                .arprot
		.hps_0_h2f_lw_axi_master_arvalid                       (hps_0_h2f_lw_axi_master_arvalid),                                //                                                .arvalid
		.hps_0_h2f_lw_axi_master_arready                       (hps_0_h2f_lw_axi_master_arready),                                //                                                .arready
		.hps_0_h2f_lw_axi_master_rid                           (hps_0_h2f_lw_axi_master_rid),                                    //                                                .rid
		.hps_0_h2f_lw_axi_master_rdata                         (hps_0_h2f_lw_axi_master_rdata),                                  //                                                .rdata
		.hps_0_h2f_lw_axi_master_rresp                         (hps_0_h2f_lw_axi_master_rresp),                                  //                                                .rresp
		.hps_0_h2f_lw_axi_master_rlast                         (hps_0_h2f_lw_axi_master_rlast),                                  //                                                .rlast
		.hps_0_h2f_lw_axi_master_rvalid                        (hps_0_h2f_lw_axi_master_rvalid),                                 //                                                .rvalid
		.hps_0_h2f_lw_axi_master_rready                        (hps_0_h2f_lw_axi_master_rready),                                 //                                                .rready
		.clock_bridge_0_out_clk_clk                            (mem_clk_clk),                                                    //                          clock_bridge_0_out_clk.clk
		.pll_reconfig_0_mgmt_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // pll_reconfig_0_mgmt_reset_reset_bridge_in_reset.reset
		.mm_bridge_h2f_lw_s0_address                           (mm_interconnect_0_mm_bridge_h2f_lw_s0_address),                  //                             mm_bridge_h2f_lw_s0.address
		.mm_bridge_h2f_lw_s0_write                             (mm_interconnect_0_mm_bridge_h2f_lw_s0_write),                    //                                                .write
		.mm_bridge_h2f_lw_s0_read                              (mm_interconnect_0_mm_bridge_h2f_lw_s0_read),                     //                                                .read
		.mm_bridge_h2f_lw_s0_readdata                          (mm_interconnect_0_mm_bridge_h2f_lw_s0_readdata),                 //                                                .readdata
		.mm_bridge_h2f_lw_s0_writedata                         (mm_interconnect_0_mm_bridge_h2f_lw_s0_writedata),                //                                                .writedata
		.mm_bridge_h2f_lw_s0_burstcount                        (mm_interconnect_0_mm_bridge_h2f_lw_s0_burstcount),               //                                                .burstcount
		.mm_bridge_h2f_lw_s0_byteenable                        (mm_interconnect_0_mm_bridge_h2f_lw_s0_byteenable),               //                                                .byteenable
		.mm_bridge_h2f_lw_s0_readdatavalid                     (mm_interconnect_0_mm_bridge_h2f_lw_s0_readdatavalid),            //                                                .readdatavalid
		.mm_bridge_h2f_lw_s0_waitrequest                       (mm_interconnect_0_mm_bridge_h2f_lw_s0_waitrequest),              //                                                .waitrequest
		.mm_bridge_h2f_lw_s0_debugaccess                       (mm_interconnect_0_mm_bridge_h2f_lw_s0_debugaccess),              //                                                .debugaccess
		.pll_reconfig_0_mgmt_avalon_slave_address              (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address),     //                pll_reconfig_0_mgmt_avalon_slave.address
		.pll_reconfig_0_mgmt_avalon_slave_write                (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write),       //                                                .write
		.pll_reconfig_0_mgmt_avalon_slave_read                 (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read),        //                                                .read
		.pll_reconfig_0_mgmt_avalon_slave_readdata             (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                                                .readdata
		.pll_reconfig_0_mgmt_avalon_slave_writedata            (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                                                .writedata
		.pll_reconfig_0_mgmt_avalon_slave_waitrequest          (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest)  //                                                .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (mem_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
